parameter M=25;
parameter N=64;
parameter K=64;
