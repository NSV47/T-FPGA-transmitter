//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.09
//Part Number: GW1NSR-LV4CQN48PC6/I5
//Device: GW1NSR-4C
//Created Time: Thu Nov 28 12:37:03 2024

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [11:0] dout;
input clk;
input oce;
input ce;
input reset;
input [11:0] ad;

wire [27:0] prom_inst_0_dout_w;
wire [27:0] prom_inst_1_dout_w;
wire [27:0] prom_inst_2_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h51EB852FB852FC962FC9630D9630DA730DA741DA741EB841EB852EB852FC852F;
defparam prom_inst_0.INIT_RAM_01 = 256'hB852FC9630C9630DA741DA741EB852EB852FC962FC9630DA630DA741EA741EB8;
defparam prom_inst_0.INIT_RAM_02 = 256'hEB852FC9630DA741EB852FC9630DA630DA741EB852FC9630C9630DA741EB851E;
defparam prom_inst_0.INIT_RAM_03 = 256'hB9630DA741EB8630DA741EB852FC9741EB852FC9630DA741EB852FC9630DA741;
defparam prom_inst_0.INIT_RAM_04 = 256'h1EC9631EB8530DA752FC9641EB8630DA752FC9631EB852FDA741EB8630DA741E;
defparam prom_inst_0.INIT_RAM_05 = 256'hEB8631EB9631EB9631EC9641EB9631EB9631EB8630EB8530DA8520DA752FC974;
defparam prom_inst_0.INIT_RAM_06 = 256'hFDA8531EC9742FDA8530EB9641FCA7520DB8631EC9641FCA752FDA8520DB8530;
defparam prom_inst_0.INIT_RAM_07 = 256'h420EB97520EC97520EC97520EC97520EB97420DB9642FDA8631FCA7530EB9642;
defparam prom_inst_0.INIT_RAM_08 = 256'hB97531FDB97531FDB97531FCA86420ECA8531FDB96420ECA7531FCA8642FDB96;
defparam prom_inst_0.INIT_RAM_09 = 256'h320ECA975320ECA975310ECA86431FDB976420ECA86431FDB97531FDB97531FD;
defparam prom_inst_0.INIT_RAM_0A = 256'hB9865320FDCA976431FECB9864310ECB986431FECA975420FDBA86531FECA875;
defparam prom_inst_0.INIT_RAM_0B = 256'h10FDCBA87653210EDCB98754310FDCB98754310FDCA9865321FECB9875421FEC;
defparam prom_inst_0.INIT_RAM_0C = 256'h543210FEDDCBA9876543210FEDCB9876543210FEDCA987654310FEDCA9876532;
defparam prom_inst_0.INIT_RAM_0D = 256'h65544322100FEEDCCBA99877654432110FEEDCBAA987665432100FEDCBA99876;
defparam prom_inst_0.INIT_RAM_0E = 256'h4433322211000FFFEEDDDCCBBBAA99887766555443221100FFEEDDCBBAA98877;
defparam prom_inst_0.INIT_RAM_0F = 256'hEEEEEEEEEEEEEEDDDDDDDDDDCCCCCCCCBBBBBBAAAAA999988887777666655544;
defparam prom_inst_0.INIT_RAM_10 = 256'h45556666777788889999AAAAABBBBBBCCCCCCCCDDDDDDDDDDEEEEEEEEEEEEEEE;
defparam prom_inst_0.INIT_RAM_11 = 256'h7889AABBCDDEEFF00112234455566778899AABBBCCDDDEEFFF00011222333444;
defparam prom_inst_0.INIT_RAM_12 = 256'h7899ABCDEF001234566789AABCDEEF01123445677899ABCCDEEF001223445567;
defparam prom_inst_0.INIT_RAM_13 = 256'h356789ACDEF013456789ACDEF0123456789BCDEF0123456789ABCDDEF0123456;
defparam prom_inst_0.INIT_RAM_14 = 256'hEF1245789BCEF1235689ACDF01345789BCDF01345789BCDE01235678ABCDF012;
defparam prom_inst_0.INIT_RAM_15 = 256'h78ACEF13568ABDF024579ACEF134689BCE0134689BCEF134679ACDF0235689BC;
defparam prom_inst_0.INIT_RAM_16 = 256'hF13579BDF13579BDF13468ACE024679BDF13468ACE013579ACE023579ACE0235;
defparam prom_inst_0.INIT_RAM_17 = 256'h9BDF2468ACF1357ACE02469BDF1358ACE02468ACF13579BDF13579BDF13579BD;
defparam prom_inst_0.INIT_RAM_18 = 256'h469BE0357ACF1368ADF2469BD02479BE02579CE02579CE02579CE02579BE0246;
defparam prom_inst_0.INIT_RAM_19 = 256'h358BD0258ADF257ACF1469CE1368BD0257ACF1469BE0358ADF2479CE1358ADF2;
defparam prom_inst_0.INIT_RAM_1A = 256'h79CF257AD0258AD0358BE0368BE1369BE1369BE1469CE1369BE1369BE1368BE0;
defparam prom_inst_0.INIT_RAM_1B = 256'h147AD0368BE147ADF258BE1369CF257AD0368BE1469CF257AD0358BE1369CE14;
defparam prom_inst_0.INIT_RAM_1C = 256'h47AD0369CF258BE147AD0369CF258BE1479CF258BE147AD0368BE147AD0369BE;
defparam prom_inst_0.INIT_RAM_1D = 256'h158BE147AD0369C0369CF258BE147AD036AD0369CF258BE147AD0369CF258BE1;
defparam prom_inst_0.INIT_RAM_1E = 256'hBE147AE147AD036AD0369CF269CF258BE258BE147AD147AD0369C0369CF258BE;
defparam prom_inst_0.INIT_RAM_1F = 256'h258CF258BE258BE148BE147AD147AD037AD0369D0369CF269CF258BF258BE158;
defparam prom_inst_0.INIT_RAM_20 = 256'h9D0369CF369CF258CF258BE158BE147BE147AD147AD036AD0369C0369CF269CF;
defparam prom_inst_0.INIT_RAM_21 = 256'h369CF258BE258BE147AD147AD0369C0369CF258CF258BE148BE147AD047AD036;
defparam prom_inst_0.INIT_RAM_22 = 256'h0369CF258BE147AD0369CF258BE148BE147AD0369CF258BE258BE147AD0369D0;
defparam prom_inst_0.INIT_RAM_23 = 256'h358BE147AD0368BE147AD0369CF257AD0369CF258BE147AD0369CF258BE147AD;
defparam prom_inst_0.INIT_RAM_24 = 256'hD0258BD0369BE1479CF258AD0368BE1479CF258BD0369CF147AD0368BE147AD0;
defparam prom_inst_0.INIT_RAM_25 = 256'h0368BD0358BD0358BD0258AD0358BD0358BD0368BE0369BE1469CE1479CF257A;
defparam prom_inst_0.INIT_RAM_26 = 256'hF1469BD0257ACF1469BE0358ADF2479CE1368BD0258ADF2479CF1469CE1369BE;
defparam prom_inst_0.INIT_RAM_27 = 256'hACE03579CE02579CE02579CE02579CE0357ACE1358ACF1468BDF2479BE0358AC;
defparam prom_inst_0.INIT_RAM_28 = 256'h3579BDF13579BDF13579BDF2468ACE02469BDF1358ACE02479BDF2468ACF1358;
defparam prom_inst_0.INIT_RAM_29 = 256'hBCE024579BCE024579BDE02468ABDF13578ACE02468ABDF13579BDF13579BDF1;
defparam prom_inst_0.INIT_RAM_2A = 256'h35689BCEF124578ABDF023568ABDE023568ABDF024579ACEF134689BDF024679;
defparam prom_inst_0.INIT_RAM_2B = 256'hDEF12346789BCDE01235679ABDEF1235679ABDEF1245689BCDF0235679ACDF02;
defparam prom_inst_0.INIT_RAM_2C = 256'h9ABCDEF01123456789ABCDEF012356789ABCDEF012456789ABDEF012456789BC;
defparam prom_inst_0.INIT_RAM_2D = 256'h899AABCCDEEF00122345567789AABCDDEF0012344567889ABCDEEF0123455678;
defparam prom_inst_0.INIT_RAM_2E = 256'hAABBBCCCDDEEEFFF00111223334455667788999AABCCDDEEFF00112334456677;
defparam prom_inst_0.INIT_RAM_2F = 256'h00000000000000111111111122222222333333444445555666677778888999AA;
defparam prom_inst_0.INIT_RAM_30 = 256'hA999888877776666555544444333333222222221111111111000000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h7665443321100FFEEDDCCBAA99988776655443332211100FFFEEEDDCCCBBBAAA;
defparam prom_inst_0.INIT_RAM_32 = 256'h765543210FEEDCBA9887654432100FEDDCBAA98776554322100FEEDCCBAA9987;
defparam prom_inst_0.INIT_RAM_33 = 256'hB987654210FEDBA987654210FEDCBA987653210FEDCBA98765432110FEDCBA98;
defparam prom_inst_0.INIT_RAM_34 = 256'h0FDCA9765320FDCB9865421FEDBA9765321FEDBA97653210EDCB98764321FEDC;
defparam prom_inst_0.INIT_RAM_35 = 256'h76420FDB986431FECA975420FDBA865320EDBA865320FDBA875421FECB986532;
defparam prom_inst_0.INIT_RAM_36 = 256'hFDB97531FDB97531FDBA86420ECA87531FDBA86420EDB975420ECB975420ECB9;
defparam prom_inst_0.INIT_RAM_37 = 256'h531FCA8642FDB97420ECA8531FDB96420ECA8642FDB97531FDB97531FDB97531;
defparam prom_inst_0.INIT_RAM_38 = 256'hA8530EB9742FDB8641FCA8531ECA7530EC97520EC97520EC97520EC97530ECA8;
defparam prom_inst_0.INIT_RAM_39 = 256'hB9631EC9641FC9742FDA8520DB8631EC9742FDA8530EB9641FCA7520DB9641FC;
defparam prom_inst_0.INIT_RAM_3A = 256'h752FC9741EC9641EB9630EB8630DB8530DB8530DA8520DB8530DB8530DB8630E;
defparam prom_inst_0.INIT_RAM_3B = 256'hDA741EB8630DA741FC9630DB852FC9741EB8630DA852FC9741EB9630DB8520DA;
defparam prom_inst_0.INIT_RAM_3C = 256'hA741EB852FC9630DA741EB852FC9630DA752FC9630DA741EB8630DA741EB8530;
defparam prom_inst_0.INIT_RAM_3D = 256'hD9630DA741EB852EB852FC9630DA741EB841EB852FC9630DA741EB852FC9630D;
defparam prom_inst_0.INIT_RAM_3E = 256'h30DA740DA741EB841EB852FC852FC9630C9630DA741DA741EB852EB852FC9630;
defparam prom_inst_0.INIT_RAM_3F = 256'hC962FC9630C9630DA630DA741DA741EB741EB851EB852FC852FC963FC9630D96;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hCCBBBBBAAAAA999998888887777766666555554444433333222221111100000F;
defparam prom_inst_1.INIT_RAM_01 = 256'h8888777777666665555544444333332222211111000000FFFFFEEEEEDDDDDCCC;
defparam prom_inst_1.INIT_RAM_02 = 256'h444443333332222211111000000FFFFFEEEEEDDDDDCCCCCCBBBBBAAAAA999998;
defparam prom_inst_1.INIT_RAM_03 = 256'h00000FFFFFEEEEEEDDDDDCCCCCBBBBBBAAAAA999999888887777766666655555;
defparam prom_inst_1.INIT_RAM_04 = 256'hCBBBBBBAAAAAA999998888887777776666655555544444333333222222111110;
defparam prom_inst_1.INIT_RAM_05 = 256'h666666555555444444333333222222111111000000FFFFFFEEEEEEDDDDDCCCCC;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000FFFFFFEEEEEEEDDDDDDCCCCCCCBBBBBBAAAAAA9999998888888777777;
defparam prom_inst_1.INIT_RAM_07 = 256'hAAA9999999888888877777776666666555555544444433333332222222111111;
defparam prom_inst_1.INIT_RAM_08 = 256'h2222221111111100000000FFFFFFFFEEEEEEEDDDDDDDDCCCCCCCBBBBBBBAAAAA;
defparam prom_inst_1.INIT_RAM_09 = 256'hAAA9999999998888888887777777766666666655555555444444443333333322;
defparam prom_inst_1.INIT_RAM_0A = 256'h00000000FFFFFFFFFFEEEEEEEEEEEDDDDDDDDDCCCCCCCCCCBBBBBBBBBAAAAAAA;
defparam prom_inst_1.INIT_RAM_0B = 256'h6655555555555554444444444443333333333332222222222211111111111000;
defparam prom_inst_1.INIT_RAM_0C = 256'hAAAAAA9999999999999999988888888888888877777777777777666666666666;
defparam prom_inst_1.INIT_RAM_0D = 256'hDDDDDDDDDDDCCCCCCCCCCCCCCCCCCCCCCBBBBBBBBBBBBBBBBBBBBAAAAAAAAAAA;
defparam prom_inst_1.INIT_RAM_0E = 256'hFFFFFFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDD;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_11 = 256'hDDDDDDDDDDDDDDDEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_12 = 256'hAAAAAAAAAABBBBBBBBBBBBBBBBBBBBCCCCCCCCCCCCCCCCCCCCCCDDDDDDDDDDDD;
defparam prom_inst_1.INIT_RAM_13 = 256'h666666666667777777777777788888888888888899999999999999999AAAAAAA;
defparam prom_inst_1.INIT_RAM_14 = 256'h0011111111111222222222223333333333334444444444445555555555555666;
defparam prom_inst_1.INIT_RAM_15 = 256'hAAAAAABBBBBBBBBCCCCCCCCCCDDDDDDDDDEEEEEEEEEEEFFFFFFFFFF000000000;
defparam prom_inst_1.INIT_RAM_16 = 256'h233333333444444445555555566666666677777777888888888999999999AAAA;
defparam prom_inst_1.INIT_RAM_17 = 256'hAAAABBBBBBBCCCCCCCDDDDDDDDEEEEEEEFFFFFFFF00000000111111112222222;
defparam prom_inst_1.INIT_RAM_18 = 256'h111112222222333333344444455555556666666777777788888889999999AAAA;
defparam prom_inst_1.INIT_RAM_19 = 256'h777778888888999999AAAAAABBBBBBCCCCCCCDDDDDDEEEEEEEFFFFFF00000001;
defparam prom_inst_1.INIT_RAM_1A = 256'hCCCCDDDDDEEEEEEFFFFFF0000001111112222223333334444445555556666667;
defparam prom_inst_1.INIT_RAM_1B = 256'h11111222222333333444445555556666677777788888899999AAAAAABBBBBBCC;
defparam prom_inst_1.INIT_RAM_1C = 256'h55556666667777788888999999AAAAABBBBBBCCCCCDDDDDEEEEEEFFFFF000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h99999AAAAABBBBBCCCCCCDDDDDEEEEEFFFFF0000001111122222333333444445;
defparam prom_inst_1.INIT_RAM_1E = 256'hCCDDDDDEEEEEFFFFF00000011111222223333344444555556666677777788888;
defparam prom_inst_1.INIT_RAM_1F = 256'h000001111122222333334444455555666667777788888899999AAAAABBBBBCCC;
defparam prom_inst_1.INIT_RAM_20 = 256'h334444445555566666777778888899999AAAAABBBBBCCCCCDDDDDEEEEEEFFFFF;
defparam prom_inst_1.INIT_RAM_21 = 256'h777778888899999AAAAABBBBBCCCCCDDDDDDEEEEEFFFFF000001111122222333;
defparam prom_inst_1.INIT_RAM_22 = 256'hBBBBBBCCCCCDDDDDEEEEEEFFFFF0000011111222222333334444455555666667;
defparam prom_inst_1.INIT_RAM_23 = 256'hFFFFF000001111112222233333344444555555666667777788888899999AAAAA;
defparam prom_inst_1.INIT_RAM_24 = 256'h344444455555566666677777888888999999AAAAABBBBBBCCCCCDDDDDDEEEEEF;
defparam prom_inst_1.INIT_RAM_25 = 256'h999999AAAAAABBBBBBCCCCCCDDDDDDEEEEEEFFFFFF0000001111112222223333;
defparam prom_inst_1.INIT_RAM_26 = 256'hEFFFFFF000000011111122222223333334444445555555666666777777888888;
defparam prom_inst_1.INIT_RAM_27 = 256'h5556666666777777788888889999999AAAAAAABBBBBBBCCCCCCCDDDDDDEEEEEE;
defparam prom_inst_1.INIT_RAM_28 = 256'hDDDDDDDEEEEEEEEFFFFFFFF00000001111111122222223333333344444445555;
defparam prom_inst_1.INIT_RAM_29 = 256'h55566666666677777777788888888899999999AAAAAAAAABBBBBBBBCCCCCCCCD;
defparam prom_inst_1.INIT_RAM_2A = 256'hFFFFFFFFF0000000000111111111122222222223333333333444444444555555;
defparam prom_inst_1.INIT_RAM_2B = 256'h999AAAAAAAAAAAABBBBBBBBBBBBBCCCCCCCCCCCCDDDDDDDDDDDEEEEEEEEEEEFF;
defparam prom_inst_1.INIT_RAM_2C = 256'h5555555666666666666666667777777777777778888888888888899999999999;
defparam prom_inst_1.INIT_RAM_2D = 256'h2222222222223333333333333333333333444444444444444444445555555555;
defparam prom_inst_1.INIT_RAM_2E = 256'h0000000000000000111111111111111111111111111111111122222222222222;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_31 = 256'h2222222222222111111111111111111111111111111111100000000000000000;
defparam prom_inst_1.INIT_RAM_32 = 256'h5555555554444444444444444444433333333333333333333332222222222222;
defparam prom_inst_1.INIT_RAM_33 = 256'h9999999999888888888888887777777777777776666666666666666655555555;
defparam prom_inst_1.INIT_RAM_34 = 256'hFEEEEEEEEEEEDDDDDDDDDDDCCCCCCCCCCCCBBBBBBBBBBBBBAAAAAAAAAAAA9999;
defparam prom_inst_1.INIT_RAM_35 = 256'h555554444444443333333333222222222211111111110000000000FFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_36 = 256'hCCCCCCCCBBBBBBBBAAAAAAAAA999999998888888887777777776666666665555;
defparam prom_inst_1.INIT_RAM_37 = 256'h5554444444333333332222222111111110000000FFFFFFFFEEEEEEEEDDDDDDDD;
defparam prom_inst_1.INIT_RAM_38 = 256'hEEEEEDDDDDDCCCCCCCBBBBBBBAAAAAAA99999998888888777777766666665555;
defparam prom_inst_1.INIT_RAM_39 = 256'h88888777777666666555555544444433333322222221111110000000FFFFFFEE;
defparam prom_inst_1.INIT_RAM_3A = 256'h333222222111111000000FFFFFFEEEEEEDDDDDDCCCCCCBBBBBBAAAAAA9999998;
defparam prom_inst_1.INIT_RAM_3B = 256'hEEEEEDDDDDDCCCCCBBBBBBAAAAA9999998888887777766666655555544444433;
defparam prom_inst_1.INIT_RAM_3C = 256'hAAAA999998888887777766666555555444443333332222211111100000FFFFFF;
defparam prom_inst_1.INIT_RAM_3D = 256'h666665555544444333332222221111100000FFFFFEEEEEEDDDDDCCCCCBBBBBBA;
defparam prom_inst_1.INIT_RAM_3E = 256'h33222221111100000FFFFFEEEEEDDDDDDCCCCCBBBBBAAAAA9999988888777777;
defparam prom_inst_1.INIT_RAM_3F = 256'hFFFFEEEEEEDDDDDCCCCCBBBBBAAAAA9999988888777776666655555444444333;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[27:0],dout[11:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 4;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h8888888888888888888888888888888888888888888888888888888888888887;
defparam prom_inst_2.INIT_RAM_01 = 256'h9999999999999999999999999999999999999999999999888888888888888888;
defparam prom_inst_2.INIT_RAM_02 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAA9999999999999999999999999999999999999;
defparam prom_inst_2.INIT_RAM_03 = 256'hBBBBBAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_2.INIT_RAM_04 = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_05 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_06 = 256'hDDDDDDDCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_07 = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD;
defparam prom_inst_2.INIT_RAM_08 = 256'hEEEEEEEEEEEEEEEEEEEEEEDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD;
defparam prom_inst_2.INIT_RAM_09 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_0A = 256'hFFFFFFFFEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_13 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_14 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_15 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_16 = 256'hEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_17 = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDEEEEEEEEEEEEEEEEEEEEEEE;
defparam prom_inst_2.INIT_RAM_18 = 256'hDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD;
defparam prom_inst_2.INIT_RAM_19 = 256'hCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCDDDDDDDD;
defparam prom_inst_2.INIT_RAM_1A = 256'hBBBBBBBBBBBBBBBBBBBBBCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC;
defparam prom_inst_2.INIT_RAM_1B = 256'hBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB;
defparam prom_inst_2.INIT_RAM_1C = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABBBBBB;
defparam prom_inst_2.INIT_RAM_1D = 256'h999999999999999999999999999999999999AAAAAAAAAAAAAAAAAAAAAAAAAAAA;
defparam prom_inst_2.INIT_RAM_1E = 256'h8888888888888888899999999999999999999999999999999999999999999999;
defparam prom_inst_2.INIT_RAM_1F = 256'h8888888888888888888888888888888888888888888888888888888888888888;
defparam prom_inst_2.INIT_RAM_20 = 256'h7777777777777777777777777777777777777777777777777777777777777777;
defparam prom_inst_2.INIT_RAM_21 = 256'h6666666666666666666666666666666666666666666666777777777777777777;
defparam prom_inst_2.INIT_RAM_22 = 256'h5555555555555555555555555556666666666666666666666666666666666666;
defparam prom_inst_2.INIT_RAM_23 = 256'h4444455555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_2.INIT_RAM_24 = 256'h4444444444444444444444444444444444444444444444444444444444444444;
defparam prom_inst_2.INIT_RAM_25 = 256'h3333333333333333333333333333333333333333334444444444444444444444;
defparam prom_inst_2.INIT_RAM_26 = 256'h2222222333333333333333333333333333333333333333333333333333333333;
defparam prom_inst_2.INIT_RAM_27 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam prom_inst_2.INIT_RAM_28 = 256'h1111111111111111111111122222222222222222222222222222222222222222;
defparam prom_inst_2.INIT_RAM_29 = 256'h1111111111111111111111111111111111111111111111111111111111111111;
defparam prom_inst_2.INIT_RAM_2A = 256'h0000000001111111111111111111111111111111111111111111111111111111;
defparam prom_inst_2.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_35 = 256'h1111111111111111111111111111111111111111111111111111110000000000;
defparam prom_inst_2.INIT_RAM_36 = 256'h1111111111111111111111111111111111111111111111111111111111111111;
defparam prom_inst_2.INIT_RAM_37 = 256'h2222222222222222222222222222222222222222111111111111111111111111;
defparam prom_inst_2.INIT_RAM_38 = 256'h2222222222222222222222222222222222222222222222222222222222222222;
defparam prom_inst_2.INIT_RAM_39 = 256'h3333333333333333333333333333333333333333333333333333333322222222;
defparam prom_inst_2.INIT_RAM_3A = 256'h4444444444444444444443333333333333333333333333333333333333333333;
defparam prom_inst_2.INIT_RAM_3B = 256'h4444444444444444444444444444444444444444444444444444444444444444;
defparam prom_inst_2.INIT_RAM_3C = 256'h5555555555555555555555555555555555555555555555555555555555444444;
defparam prom_inst_2.INIT_RAM_3D = 256'h6666666666666666666666666666666666665555555555555555555555555555;
defparam prom_inst_2.INIT_RAM_3E = 256'h7777777777777777766666666666666666666666666666666666666666666666;
defparam prom_inst_2.INIT_RAM_3F = 256'h7777777777777777777777777777777777777777777777777777777777777777;

endmodule //Gowin_pROM
